`timescale 1ns / 1ns		//仿真时间单位/时间精度
module testbench();		//信号声明
	reg f0,clk;
	wire f1;
	
	parameter T = 20;	//初始周期20ns
	initial		//复位
	begin
		clk = 0;
	end
	initial
	begin//25组f0
		f0=0;
		#10000
		f0=1;
		#40000
		f0=0;
		#15000
		f0=1;
		#35000
		f0=0;
		#20000
		f0=1;
		#30000
		f0=0;
		#30000
		f0=1;
		#20000
		f0=0;
		#25000
		f0=1;
		#25000
		f0=0;
		#10000
		f0=1;
		#40000
		f0=0;
		#15000
		f0=1;
		#35000
		f0=0;
		#20000
		f0=1;
		#30000
		f0=0;
		#30000
		f0=1;
		#20000
		f0=0;
		#25000
		f0=1;
		#25000
		f0=0;
		#10000
		f0=1;
		#40000
		f0=0;
		#15000
		f0=1;
		#35000
		f0=0;
		#20000
		f0=1;
		#30000
		f0=0;
		#30000
		f0=1;
		#20000
		f0=0;
		#25000
		f0=1;
		#25000
		f0=0;
		#10000
		f0=1;
		#40000
		f0=0;
		#15000
		f0=1;
		#35000
		f0=0;
		#20000
		f0=1;
		#30000
		f0=0;
		#30000
		f0=1;
		#20000
		f0=0;
		#25000
		f0=1;
		#25000
		f0=0;
		#10000
		f0=1;
		#40000
		f0=0;
		#15000
		f0=1;
		#35000
		f0=0;
		#20000
		f0=1;
		#30000
		f0=0;
		#30000
		f0=1;
		#20000
		f0=0;
		#25000
		f0=1;
		//#25000
	end
	always #(T/2)
		clk=~clk;
	dcl_1778_6 divider(
		.clk(clk),
		.f0(f0),
		.f1(f1)
	);
endmodule